module Arithmetic(X,Y, sel, out);
input [3:0] X,Y;
input [1:0] sel;
output [7:0] out;

reg tempOut;

assign out = 5;

endmodule 